$date
	Tue Oct 14 18:58:46 2025
$end
$version
	Icarus Verilog
$end
$timescale
	1ns
$end
$scope module decoder_2_4_tb $end
$var wire 4 ! y [3:0] $end
$var reg 2 " I [1:0] $end
$var reg 1 # e $end
$scope module decoder_2_4_1 $end
$var wire 2 $ I [1:0] $end
$var wire 1 # e $end
$var reg 4 % y [3:0] $end
$upscope $end
$upscope $end
$enddefinitions $end
$comment Show the parameter values. $end
$dumpall
$end
#0
$dumpvars
b1 %
b0 $
1#
b0 "
b1 !
$end
#10
b10 !
b10 %
b1 "
b1 $
#20
b100 !
b100 %
b10 "
b10 $
#30
b1000 !
b1000 %
b11 "
b11 $
#40
b0 !
b0 %
b0 "
b0 $
0#
#50
